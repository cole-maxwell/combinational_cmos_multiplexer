    Mac OS X            	   2   �      �                                      ATTR       �   �   H                  �   H  com.apple.macl    ����&�H��Y/ 24O� �hg�D����#�:CU                                    