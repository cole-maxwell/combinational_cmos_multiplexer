* First line is treated as comment
.options list node post
* Include transistor models. include command can also be used to include other spice files
.include '$PDK_DIR/ncsu_basekit/models/hspice/hspice_nom.include'

.param vdd_val=0.8

Vsupply vdd 0 vdd_val
Vgnd GND 0 0

* Digital vector file for input
.vec 'input.vec'

.subckt inverter GND VDD IN OUT size=1
m0 out in vdd vdd PMOS_VTL L=50e-9 W='size*180e-9'
m1 out in 0   0   NMOS_VTL L=50e-9 W='size*90e-9'
.ends


Xinv_1 GND VDD A A_bar inverter size=1
Xinv_2 GND VDD B B_bar inverter size=1.5


Cload B_bar 0 1e-15

.tran 1p 0.5n

* .measure can be used for power, delay measurements

.end
